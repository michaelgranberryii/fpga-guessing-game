`timescale 1ns / 1ps
module debounce_tb;
    
endmodule
