module single_pulse_detector_tb;

endmodule